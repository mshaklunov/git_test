
module

always @(posedge clk)
begin

counter<= counter+1;

end

endmodule
